`include "logical/rtl/axi4_lite_master.v"
`include "logical/rtl/axi4_lite_slave.v"
`include "logical/rtl/axi4_lite_interconnect/axi4_lite_interconnect_m1s2.v"
`include "logical/rtl/wrapper/axi4_lite_master_wrapper.v"
`include "logical/rtl/wrapper/axi4_lite_slave_wrapper.v"
`include "logical/tb/tb_wrapper/dummy/handler/master.v"
`include "logical/tb/tb_wrapper/dummy/handler/slave.v"
`include "logical/tb/tb_wrapper/dummy/wrapper/dut_axi4_lite_master_wrapper.v"
`include "logical/tb/tb_wrapper/dummy/wrapper/dut_axi4_lite_slave_wrapper.v"
// `include "logical/tb/tb_wrapper/tb_wrapper_master.v"
// `include "logical/tb/tb_wrapper/tb_wrapper_slave.v"
